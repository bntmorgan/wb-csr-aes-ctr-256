`define AES_CSR_CTRL 10'h000
`define AES_CSR_STAT 10'h001
`define AES_CSR_KEY0 10'h010
`define AES_CSR_KEY1 10'h011
`define AES_CSR_KEY2 10'h012
`define AES_CSR_KEY3 10'h013
`define AES_CSR_KEY4 10'h014
`define AES_CSR_KEY5 10'h015
`define AES_CSR_KEY6 10'h016
`define AES_CSR_KEY7 10'h017
`define AES_CSR_NONC 10'h021
`define AES_CSR_IV_0 10'h022
`define AES_CSR_IV_1 10'h023

`define AES_STATE_IDLE 1'b0
`define AES_STATE_RUN  1'b1
